module dht11_function (
    ports
);
    
endmodule

