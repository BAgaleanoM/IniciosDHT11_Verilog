module DataReciverModule (
    input wire clk,
    input wire rst,
    input reg[39:0] data_dht11, //Variable que almacena la cadena de bits, luego de las señales de checkeo
    output reg[15:0] temp_data,
    output reg[15:0] hum_data
);



endmodule
