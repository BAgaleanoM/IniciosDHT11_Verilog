module moduleName (
    input wire clk,
    input wire rst,

);



endmodule
