
module StartModule (
    input wire clk,
    input wire rst,
    input wire 
);
    
endmodule